`include "../../common/hdl/bcpu_cond_defs.vh"


`define ALUOP_ADDNF    4'b0000
`define ALUOP_SUBNF    4'b0001
`define ALUOP_ADD      4'b0010
`define ALUOP_ADC      4'b0011
`define ALUOP_SUB      4'b0100
`define ALUOP_SBC      4'b0101
`define ALUOP_RSUB     4'b0110
`define ALUOP_RSBC     4'b0111
`define ALUOP_AND      4'b1000
`define ALUOP_ANDN     4'b1001
`define ALUOP_OR       4'b1010
`define ALUOP_XOR      4'b1011
`define ALUOP_MUL      4'b1100
`define ALUOP_MULHSU   4'b1101
`define ALUOP_MULHUU   4'b1110
`define ALUOP_MULHSS   4'b1111


