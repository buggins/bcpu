`include "../../common/hdl/bcpu_cond_defs.vh"

`define MUL_B_SIGN 3
`define MUL_A_SIGN 2

`define ALUOP_INC  4'b0000
`define ALUOP_DEC  4'b0001
`define ALUOP_ADD  4'b0010
`define ALUOP_ADC  4'b0011
`define ALUOP_SUB  4'b0100
`define ALUOP_SBC  4'b0101
`define ALUOP_RSUB 4'b0110
`define ALUOP_RSBC 4'b0111
`define ALUOP_AND  4'b1000
`define ALUOP_ANDN 4'b1001
`define ALUOP_OR   4'b1010
`define ALUOP_XOR  4'b1011
`define ALUOP_RES0 4'b1100
`define ALUOP_RES1 4'b1101
`define ALUOP_RES2 4'b1110
`define ALUOP_RES3 4'b1111

